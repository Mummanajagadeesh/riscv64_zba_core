//------------------------------------------------------------------------------
// File Name  : result_mux.sv
// Author     : Jagadeesh Mummana
// Email      : mummanajagadeesh97@gmail.com
// Repository : Mummanajagadeesh /riscv64_zba_core
//
// Description:
// This module implements the write-back result selection multiplexer.
// It selects the final value to be written to the register file based
// on the result source control signal.
//
// Key Features:
// - Supports ALU result write-back
// - Supports load data write-back
// - Supports PC+4 write-back for control-flow instructions
// - Supports immediate-based write-back
//
// Assumptions & Notes:
// - ResultSrcW encoding is generated by the control logic
// - Only one result source is selected per instruction
//------------------------------------------------------------------------------


module result_mux (
    input  [63:0] ALUResultW,   // ALU result (write-back stage)
    input  [63:0] ReadDataW,    // Memory read data (write-back stage)
    input  [63:0] PCPlus4W,     // PC + 4 (write-back stage)
    input  [63:0] ExtImmW,      // Immediate value (write-back stage)
    input  [1:0]  ResultSrcW,   // Result source select
    output [63:0] ResultW       // Selected write-back result
);

  // --------------------------------------------------
  // Write-back result selection
  // --------------------------------------------------
  // Selects the appropriate result based on the control
  // signal provided by the decode logic.
  assign ResultW =
      (ResultSrcW == 2'b00) ? ALUResultW :
      (ResultSrcW == 2'b01) ? ReadDataW  :
      (ResultSrcW == 2'b10) ? PCPlus4W   :
                              ExtImmW;

endmodule


//------------------------------------------------------------------------------
// Functional Summary:
// This result multiplexer determines the final value written to the register
// file, enabling correct completion of arithmetic, memory, control-flow,
// and immediate-based instructions.
//------------------------------------------------------------------------------
