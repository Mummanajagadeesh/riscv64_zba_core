//------------------------------------------------------------------------------
// File Name  : mux_SrcAE.sv
// Author     : Jagadeesh Mummana
// Email      : mummanajagadeesh97@gmail.com
// Repository : Mummanajagadeesh /riscv64_zba_core
//
// Description:
// This module implements the forwarding multiplexer for the ALU source A
// operand in the execute stage. It selects the appropriate operand based on
// forwarding control signals to resolve data hazards.
//
// Key Features:
// - Supports forwarding from MEM and WB pipeline stages
// - Combinational selection logic
// - Prevents pipeline stalls for most data hazards
//
// Assumptions & Notes:
// - ForwardAE encoding is generated by the hazard unit
// - Default selection uses register file output
//------------------------------------------------------------------------------


module mux_SrcAE (
    input  [63:0] RD1E,        // Register file source operand (execute stage)
    input  [63:0] ResultW,     // Write-back stage result
    input  [63:0] ALUResultM,  // Memory stage ALU result
    input  [1:0]  ForwardAE,   // Forwarding select control
    output [63:0] SrcAE        // Selected ALU source A
);

  // --------------------------------------------------
  // Forwarding multiplexer logic
  // --------------------------------------------------
  // Selects the correct source operand based on the
  // forwarding control encoding.
  assign SrcAE =
      (ForwardAE == 2'b00) ? RD1E :       // No forwarding
      (ForwardAE == 2'b01) ? ResultW :    // Forward from WB stage
                             ALUResultM; // Forward from MEM stage

endmodule


//------------------------------------------------------------------------------
// Functional Summary:
// This forwarding multiplexer resolves execute-stage data hazards by selecting
// the most recent version of a source operand from either the register file,
// memory stage, or write-back stage.
//------------------------------------------------------------------------------
