//------------------------------------------------------------------------------
// File Name  : mux_SrcBE2.sv
// Author     : Jagadeesh Mummana
// Email      : mummanajagadeesh97@gmail.com
// Repository : Mummanajagadeesh /riscv64_zba_core
//
// Description:
// This module implements the second-stage multiplexer for ALU source B.
// It selects between a forwarded register value and an immediate operand
// based on the ALU source control signal.
//
// Key Features:
// - Supports register and immediate-based ALU operations
// - Simple combinational selection logic
// - Used in execute stage operand selection
//
// Assumptions & Notes:
// - ALUSrcE is generated by the decode/control logic
// - Immediate value is already sign-extended
//------------------------------------------------------------------------------


module mux_SrcBE2 (
    input  [63:0] WriteDataE,   // Forwarded or register-based operand
    input  [63:0] ExtImmE,       // Sign-extended immediate value
    input         ALUSrcE,       // ALU source select control
    output [63:0] SrcBE          // Selected ALU source B
);

  // --------------------------------------------------
  // ALU source B selection
  // --------------------------------------------------
  // Chooses between register-based data and immediate
  // value for ALU operations.
  assign SrcBE = ALUSrcE ? ExtImmE : WriteDataE;

endmodule


//------------------------------------------------------------------------------
// Functional Summary:
// This multiplexer selects the appropriate second operand for the ALU,
// enabling both register-register and register-immediate instruction
// execution in the execute stage.
//------------------------------------------------------------------------------
