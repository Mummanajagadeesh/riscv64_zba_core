//------------------------------------------------------------------------------
// File Name  : mux_SrcBE1.sv
// Author     : Jagadeesh Mummana
// Email      : mummanajagadeesh97@gmail.com
// Repository : Mummanajagadeesh /riscv64_zba_core
//
// Description:
// This module implements the forwarding multiplexer for the ALU source B
// operand prior to immediate selection. It selects the appropriate register
// or forwarded value to be used as write data or ALU operand.
//
// Key Features:
// - Supports forwarding from MEM and WB pipeline stages
// - Combinational selection logic
// - Used in both ALU operations and store data path
//
// Assumptions & Notes:
// - ForwardBE encoding is generated by the hazard unit
// - Default path uses register file output
//------------------------------------------------------------------------------


module mux_SrcBE1 (
    input  [63:0] RD2E,        // Register file source operand (execute stage)
    input  [63:0] ResultW,     // Write-back stage result
    input  [63:0] ALUResultM,  // Memory stage ALU result
    input  [1:0]  ForwardBE,   // Forwarding select control
    output [63:0] WriteDataE   // Selected operand before ALUSrc mux
);

  // --------------------------------------------------
  // Forwarding multiplexer logic
  // --------------------------------------------------
  // Selects the correct operand based on the forwarding
  // control encoding.
  assign WriteDataE =
      (ForwardBE == 2'b00) ? RD2E :        // No forwarding
      (ForwardBE == 2'b01) ? ResultW :     // Forward from WB stage
                             ALUResultM;  // Forward from MEM stage

endmodule


//------------------------------------------------------------------------------
// Functional Summary:
// This module resolves data hazards for the second ALU operand by forwarding
// the most recent value from later pipeline stages, ensuring correct execution
// without unnecessary pipeline stalls.
//------------------------------------------------------------------------------
