//------------------------------------------------------------------------------
// File Name  : WD3_mux.sv
// Author     : Jagadeesh Mummana
// Email      : mummanajagadeesh97@gmail.com
// Repository : Mummanajagadeesh /riscv64_zba_core
//
// Description:
// This module implements a write-back data selection multiplexer used in the
// decode stage. It selects between the sequential PC value and the computed
// execution result based on the write-back source control signal.
//
// Key Features:
// - Selects PC+4 for control-flow instructions
// - Selects execution result for regular instructions
// - Simple combinational multiplexer
//
// Assumptions & Notes:
// - WD3_SrcD is generated by the control unit
// - PCPlus4D corresponds to the decode-stage PC increment
//------------------------------------------------------------------------------


module WD3_mux (
    input [31:0] PCPlus4D,     // PC + 4 value (decode stage)
    ResultW,                    // Execution result value
    input WD3_SrcD,             // Write-back source select
    output [31:0] OUTWD3        // Selected write-back data
);

  // --------------------------------------------------
  // Write-back data selection
  // --------------------------------------------------
  // Selects between PC+4 and execution result based
  // on the control signal.
  assign OUTWD3 = WD3_SrcD ? PCPlus4D : ResultW;

endmodule


//------------------------------------------------------------------------------
// Functional Summary:
// This multiplexer determines the data forwarded toward the register file
// write-back path in the decode stage, enabling correct handling of
// control-flow instructions that require PC-based write-back.
//------------------------------------------------------------------------------
